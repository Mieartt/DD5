library ieee;
use.ieee_std_logic_1164.all;
entity youcef is
    port (
        KHCHAM : in std_logic;
        FOM    : out std_logic
    );
architecture chbab_YOUCEF of youcef is
signal nice_hair : std_logic;
signal head : std_logic;
begin
end chbab_YOUCEF;
