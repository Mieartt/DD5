library ieee;
use.ieee_std_logic_1164.all;
entity youcef is
    port (
        wednin : in std_logic;
        fom : out std_logic
    );
architecture chbab of youcef is
signal nice_hair : std_logic;
signal head : std_logic;
begin
end chbab;
